-- megafunction wizard: %RAM: 2-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: frame_buffer.vhd
-- Megafunction Name(s):
-- 			altsyncram
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 10.0 Build 262 08/18/2010 SP 1 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2010 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY frame_buffer IS
	PORT
	(
		data		 : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		rdaddress : IN STD_LOGIC_VECTOR (16 DOWNTO 0);
		rdclock	 : IN STD_LOGIC ;
		wraddress : IN STD_LOGIC_VECTOR (16 DOWNTO 0);
		wrclock	 : IN STD_LOGIC;
		wren		 : IN STD_LOGIC;
		q		    : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
END frame_buffer;

ARCHITECTURE SYN OF frame_buffer IS
	COMPONENT spartan_frame_buffer
	  PORT (
		 clka : IN STD_LOGIC;
		 wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
		 addra : IN STD_LOGIC_VECTOR(16 DOWNTO 0);
		 dina : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 clkb : IN STD_LOGIC;
		 addrb : IN STD_LOGIC_VECTOR(16 DOWNTO 0);
		 doutb : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	  );
	END COMPONENT;

   signal wren_vector : STD_LOGIC_VECTOR (0 DOWNTO 0);
BEGIN
   wren_vector(0)  <= wren;

fb : spartan_frame_buffer
	  PORT MAP (
		 clka => wrclock,
		 wea => wren_vector,
		 addra => wraddress,
		 dina => data,
		 clkb => rdclock,
		 addrb => rdaddress,
		 doutb => q
	  );
END SYN;
